module led(
    input [7:0] LED_in,
    output [7:0] LED_out
);

    assign LED_out = LED_in;

endmodule